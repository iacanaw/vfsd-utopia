`ifndef AGENT__UVM
`define AGENT__UVM


`endif